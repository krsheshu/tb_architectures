//-----------------------------------------------------------------------------------------------------
// Copyright: Free
// Author: krsheshu
// Brief: BFM for clk_reset
//-----------------------------------------------------------------------------------------------------


interface clk_reset_bfm

  //-------------------------------------------------------------
  //  Imports
  //-------------------------------------------------------------
  import        clock_period_pkg ::  CLKPERIOD_NS       ;

  //-------------------------------------------------------------
  //  Interface signals
  //-------------------------------------------------------------

  clk_reset_interface           clk_rst_if

  //-------------------------------------------------------------
  //  Clk Description
  //-------------------------------------------------------------

  initial begin
      clk_rst_if.clk_i   =   0;
      forever begin
        # (CLKPERIOD_NS/2);
        clk_rst_if.clk_i = ~clk_rst_if.clk_i;
      end
  end


  //-------------------------------------------------------------
  //  Initialize module input signals
  //-------------------------------------------------------------

  initial begin
      clk_rst_if.reset_n_i     =   1'b1    ;
      clk_rst_if.start_i       =   1'b0    ;
  end

  //----------------------------------------------------------------------------------
  // Task: assert reset
  //----------------------------------------------------------------------------------

  task assert_reset ( )

      clk_rst_if.reset_n_i     =   1'b0    ;

  endtask : assert_reset


  //----------------------------------------------------------------------------------
  // Task: deassert reset
  //----------------------------------------------------------------------------------

  task deassert_reset ( )

      clk_rst_if.reset_n_i     =   1'b1    ;

  endtask : deassert_reset

  //----------------------------------------------------------------------------------
  // Task: assert_reset_clks
  //----------------------------------------------------------------------------------

  task assert_reset_clks ( integer nb_clks )

      assert_reset ();
      repeat ( nb_clks ) @ ( posedge clk_rst_if.clk_i );
      deassert_reset ();

  endtask : reset_module

//----------------------------------------------------------------------------------
endinterface : clk_reset_bfm
