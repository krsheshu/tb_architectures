//-----------------------------------------------------------------------------------------------------
// Copyright: Free
// Author: krsheshu
// Brief: tiny_alu_interface
//-----------------------------------------------------------------------------------------------------

interface clk_reset_interface

  //-------------------------------------------------------------
  //  Interface Signals
  //-------------------------------------------------------------

  logic                            clk_i        ;
  logic                            reset_n_i    ;

//-----------------------------------------------------------------------------------------------------

endinterface : clk_reset_interface

//-----------------------------------------------------------------------------------------------------
