//-----------------------------------------------------------------------------------------------------
// Copyright: Free
// Author: krsheshu
// Brief: BFM for tiny_alu
//-----------------------------------------------------------------------------------------------------


interface tiny_alu_bfm

  //-------------------------------------------------------------
  //  Imports
  //-------------------------------------------------------------
  import        clock_period_pkg ::  CLKPERIOD_NS             ;

  //-------------------------------------------------------------
  //  Ports
  //-------------------------------------------------------------
  (
      input   logic                            clk_i        ;
      input   logic                            reset_n_i
  );
  //-------------------------------------------------------------
  //  Interface signals
  //-------------------------------------------------------------
   (

      tiny_alu_intf         intf

   );

  //-------------------------------------------------------------
  //  Clk Description
  //-------------------------------------------------------------

  initial begin
      intf.clk_i   =   0;
      forever begin
        # (CLKPERIOD_NS/2);
        intf.clk_i = ~intf.clk_i;
      end
  end


  //-------------------------------------------------------------
  //  Initialize module input signals
  //-------------------------------------------------------------

  initial begin
      intf.reset_n_i     =   1'b1    ;
      intf.start_i       =   1'b0    ;
  end

  //----------------------------------------------------------------------------------
  // Task: assert reset
  //----------------------------------------------------------------------------------

  task assert_reset ( integer nb_clks )

      intf.reset_n_i     =   1'b0    ;
      intf.reset_n_i     =   repeat ( nb_clks ) @posedge ( intf.clk_i ) 1'b1 ;

  endtask


  //----------------------------------------------------------------------------------
  // Task: assert reset
  //----------------------------------------------------------------------------------

  task assert_reset ( integer nb_clks )

      intf.reset_n_i     =   1'b0    ;
      intf.reset_n_i     =   repeat ( nb_clks ) @posedge ( intf.clk_i ) 1'b1 ;

  endtask






//----------------------------------------------------------------------------------
endinterface : tiny_alu_bfm
