//-----------------------------------------------------------------------------------------------------
// Copyright: Free
// Author: krsheshu
// Brief: tiny_alu_bus_interface
//-----------------------------------------------------------------------------------------------------

interface tiny_alu_bus_interface

  //-------------------------------------------------------------
  //  Imports
  //-------------------------------------------------------------

  import tiny_alu_pkg ::  OPCODE_BITS  ;

  parameter   ( INPUT_DATA_BITS     =     8   );

  //-------------------------------------------------------------
  //  Interface signals
  //-------------------------------------------------------------

  logic        [ INPUT_DATA_BITS-1: 0 ]        a_i          ;
  logic        [ INPUT_DATA_BITS-1: 0 ]        b_i          ;

  logic        [ OPCODE_BITS-1: 0 ]            opcode_i     ;
  logic                                        start_i      ;

  logic        [ INPUT_DATA_BITS*2-1: 0 ]      result_o     ;
  logic                                        done_o       ;

//-----------------------------------------------------------------------------------------------------

endinterface : tiny_alu_bus_interface

//-----------------------------------------------------------------------------------------------------
